library verilog;
use verilog.vl_types.all;
entity Output_Ports_vlg_vec_tst is
end Output_Ports_vlg_vec_tst;
